library verilog;
use verilog.vl_types.all;
entity DSP_FPGA_IMC_PMSM_vlg_vec_tst is
end DSP_FPGA_IMC_PMSM_vlg_vec_tst;
