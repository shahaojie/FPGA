module Control_CLK(
				clk_ts,		// output: h0FC01
		
				clk,			// input:clock
				global_rst	// input:global_rst		
				);
				
output clk_ts;

input clk;
input global_rst;				
				
always @ (posedge clk or negedge global_rst)				
begin
	if (!global_rst)
	begin
	
	
	
	
	
	
	
	
	end
	else
	begin
	
	
	
	
	
		
	
	end







end


				
endmodule